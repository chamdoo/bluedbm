// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemServer::*;
import MemTypes::*;
import XbsvXilinxCells::*;
import HostInterface::*;

// generated by tool
import FlashEmuRequestWrapper::*;
import PlatformRequestWrapper::*;
import DmaConfigWrapper::*;
import FlashEmuIndicationProxy::*;
import DmaIndicationProxy::*;
import PlatformIndicationProxy::*;

// defined by user
import FlashEmu::*;
import BlueDBMPlatform::*;
import PlatformInterfaces::*;
import DRAMController::*;

import Clocks          :: *;
import DefaultValue    :: *;
import XilinxVC707DDR3::*;
import Xilinx       :: *;
import XilinxCells :: *;

import AuroraImportVC707::*;
import AuroraImportVC707_625::*;
import I2CSimple::*;

typedef enum {FlashEmuIndication, FlashEmuRequest, DmaIndication, DmaConfig, PlatformIndication, PlatformRequest} IfcNames deriving (Eq,Bits);

interface BlueDBMTopPins;
	interface DDR3_Pins_VC707 ddr3;
	interface Aurora_Pins_VC707 aurora0;
	interface Aurora_Pins_VC707 aurora1_0;
	interface I2C_Pins i2c;
	method Action gtx_clk_0_p(Bit#(1) v);
	method Action gtx_clk_0_n(Bit#(1) v);
	method Action gtx_clk_1_0_p(Bit#(1) v);
	method Action gtx_clk_1_0_n(Bit#(1) v);
	interface Clock deleteme_unused_clock;
	interface Reset deleteme_unused_reset;
endinterface

interface TopParam;
   interface Clock sys_clk_200mhz;
   interface Reset pci_sys_reset_n;
endinterface

module mkTopParam#(Clock asys_clk_200mhz, Reset apci_sys_reset_n)(TopParam);
   interface Clock sys_clk_200mhz = asys_clk_200mhz;
   interface Reset pci_sys_reset_n = apci_sys_reset_n;
endmodule

typedef 1 NumMasters;
module mkPortalTop#(HostType host) (PortalTop#(addrWidth, 64, BlueDBMTopPins, NumMasters)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   PlatformIndicationProxy platformIndicationProxy <- mkPlatformIndicationProxy(PlatformIndication);
   FlashEmuIndicationProxy interfaceIndicationProxy <- mkFlashEmuIndicationProxy(FlashEmuIndication);
   FlashEmu flashEmu <- mkFlashEmu(interfaceIndicationProxy.ifc, platformIndicationProxy.ifc);
   FlashEmuRequestWrapper interfaceRequestWrapper <- mkFlashEmuRequestWrapper(FlashEmuRequest,flashEmu.request);
	

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   Vector#(NumMasters, ObjectReadClient#(64))   readClients = cons(flashEmu.dmaReadClient, nil);
   Vector#(NumMasters, ObjectWriteClient#(64)) writeClients = cons(flashEmu.dmaWriteClient, nil);
   MemServer#(addrWidth, 64, NumMasters)   dma <- mkMemServer(dmaIndicationProxy.ifc, readClients, writeClients);
   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);


`ifdef BSIM
   DRAMControllerIfc dramController <- mkDRAMControllerBSIM;
   Vector#(I2C_Count,I2C_User) i2c = ?;
`else
   //////////////// test DDR3 stuff start //////////////
   //Clock sys_clk <- mkClockIBUFDS(sys_clk_200mhz, sys_reset_200mhz);

   Vector#(AuroraPorts,Clock) gtx_clk_p;
   Vector#(AuroraPorts,Clock) gtx_clk_n;
   Vector#(AuroraPorts, B2C1) pclk;
   Vector#(AuroraPorts, B2C1) nclk;
   for(Integer i = 0; i < valueOf(AuroraPorts); i=i+1) begin
       pclk[i] <- mkB2C1();
       gtx_clk_p[i] = pclk[i].c;
       nclk[i] <- mkB2C1();
       gtx_clk_n[i] = nclk[i].c;
   end
   
   Clock defaultClock <- exposeCurrentClock();
   Reset defaultReset <- exposeCurrentReset();
   Clock sys_clk = host.tsys_clk_200mhz;
   Reset pci_sys_reset_n = host.tpci_sys_reset_n;

   ClockGenerator7Params clk_params = defaultValue();
   clk_params.clkin1_period     = 5.000;       // 200 MHz reference
   clk_params.clkin_buffer      = False;       // necessary buffer is instanced above
   clk_params.reset_stages      = 0;           // no sync on reset so input clock has pll as only load
   clk_params.clkfbout_mult_f   = 5.000;       // 1000 MHz VCO
   clk_params.clkout0_divide_f  = 10;          // unused clock 
   //clk_params.clkout0_divide_f  = 8;//10;          // unused clock 
   clk_params.clkout1_divide    = 5;           // ddr3 reference clock (200 MHz)

   ClockGenerator7 clk_gen <- mkClockGenerator7(clk_params, clocked_by sys_clk, reset_by pci_sys_reset_n);
   Clock ddr_clk = clk_gen.clkout0;
   Reset rst_n <- mkAsyncReset( 4, pci_sys_reset_n, ddr_clk );
   Reset ddr3ref_rst_n <- mkAsyncReset( 4, rst_n, clk_gen.clkout1 );
   //Reset ddr3ref_rst_n <- mkAsyncReset( 1, pci_sys_reset_n, clk_gen.clkout1 );

   DDR3_Configure ddr3_cfg = defaultValue;
   //ddr3_cfg.reads_in_flight = 2;   // adjust as needed
   ddr3_cfg.reads_in_flight = 24;   // adjust as needed
   //ddr3_cfg.fast_train_sim_only = False; // adjust if simulating
   DDR3_Controller_VC707 ddr3_ctrl <- mkDDR3Controller_VC707(ddr3_cfg, clk_gen.clkout1, clocked_by clk_gen.clkout1, reset_by ddr3ref_rst_n);

   // ddr3_ctrl.user needs to connect to user logic and should use ddr3clk and ddr3rstn
   Clock ddr3clk = ddr3_ctrl.user.clock;
   Reset ddr3rstn = ddr3_ctrl.user.reset_n;
   DRAMControllerIfc dramController <- mkDRAMController(ddr3_ctrl.user, clocked_by ddr_clk, reset_by rst_n);
   
   ///////////////////////////// DDR3 end

	Clock cur_clk <- exposeCurrentClock;
	Reset cur_rst_n <- exposeCurrentReset;

	//////////////////////////// Aurora Start
	MakeResetIfc auroraRst <- mkReset(1, False, cur_clk);
	Reset auroraRstE <- mkResetEither(auroraRst.new_rst, cur_rst_n);
	Vector#(AuroraPorts, Clock) gtx_clks;
	gtx_clks[0] <- mkClockIBUFDS_GTE2(True, gtx_clk_p[0], gtx_clk_n[0]);
	gtx_clks[1] <- mkClockIBUFDS_GTE2(True, gtx_clk_p[1], gtx_clk_n[1]);

/* jca -- remove Aurora
	Vector#(AuroraPorts, AuroraIfc) auroras;
	Aurora_V7 auroraImport0 <- mkAuroraWrapper(gtx_clks[0], cur_clk, auroraRstE);//cur_rst_n);
	AuroraIfc aurora0 <- mkAurora(auroraImport0, auroraRst);
	auroras[0] = aurora0;
	
	Aurora_V7 auroraImport1_0 <- mkAuroraWrapper625(gtx_clks[1], cur_clk, auroraRstE);//cur_rst_n);
	AuroraIfc aurora1_0 <- mkAurora(auroraImport1_0, auroraRst);
	auroras[1] = aurora1_0;
*/

	//////////////////////////// Aurora End
   
   /////FIXME: Change it to use BSV's vanilla distributed I2C
   Vector#(I2C_Count,I2C_User) i2c;
   I2C i2c0 <- mkI2C(416); //125/417 = 299khz/3 = 100khz i2c clk
   i2c[0] = i2c0.user;
   
`endif
   
   BlueDBMPlatformIfc bluedbm <- mkBlueDBMPlatform(flashEmu.flash, flashEmu.host, dramController, /*auroras,*/ i2c);
   PlatformRequestWrapper platformRequestWrapper <- mkPlatformRequestWrapper(PlatformRequest, bluedbm.request);
   
   Vector#(6,StdPortal) portals;
   portals[1] = interfaceRequestWrapper.portalIfc;
   portals[0] = interfaceIndicationProxy.portalIfc; 
   portals[3] = dmaRequestWrapper.portalIfc;
   portals[2] = dmaIndicationProxy.portalIfc; 
   portals[5] = platformRequestWrapper.portalIfc;
   portals[4] = platformIndicationProxy.portalIfc;
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   //let interrupt_mux <- mkInterruptMux(portals);

   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;


`ifndef BSIM
   //interface DDR3_Pins_VC707 pins = ddr3_ctrl.ddr3;
   interface BlueDBMTopPins pins;
	   interface DDR3_Pins_VC707 ddr3 = ddr3_ctrl.ddr3;
/* remove aurora
	   interface Aurora_Pins_VC707 aurora0 = auroraImport0.aurora;
	   interface Aurora_Pins_VC707 aurora1_0 = auroraImport1_0.aurora;
*/

	   interface I2C_Pins i2c = i2c0.i2c;
	   method Action gtx_clk_0_p(Bit#(1) v);
	      pclk[0].inputclock(v);
           endmethod
	   method Action gtx_clk_0_n(Bit#(1) v);
	      nclk[0].inputclock(v);
           endmethod
	   method Action gtx_clk_1_0_p(Bit#(1) v);
	      pclk[1].inputclock(v);
           endmethod
	   method Action gtx_clk_1_0_n(Bit#(1) v);
	      nclk[1].inputclock(v);
           endmethod
	   interface deleteme_unused_clock = defaultClock;
	   interface deleteme_unused_reset = defaultReset;
   endinterface
`endif

endmodule
